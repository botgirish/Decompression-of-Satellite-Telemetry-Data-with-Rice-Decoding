module pencoder (
    input  [63:0] in,
    input reset,
    input peen,
    output reg [9:0] out,  // Now 10-bit wide
    output reg [5:0] len   // Remains 6-bit
);

always @(*) begin
    if (reset) begin
        out <= 10'd0;
        len <= 6'd0;
    end
    else if (peen) begin
        casex (in)
            64'b1???????????????????????????????????????????????????????????????: begin out = 10'd0;  len = 6'd1;  end
            64'b01??????????????????????????????????????????????????????????????: begin out = 10'd1;  len = 6'd2;  end
            64'b001?????????????????????????????????????????????????????????????: begin out = 10'd2;  len = 6'd3;  end
            64'b0001????????????????????????????????????????????????????????????: begin out = 10'd3;  len = 6'd4;  end
            64'b00001???????????????????????????????????????????????????????????: begin out = 10'd4;  len = 6'd5;  end
            64'b000001??????????????????????????????????????????????????????????: begin out = 10'd5;  len = 6'd6;  end
            64'b0000001?????????????????????????????????????????????????????????: begin out = 10'd6;  len = 6'd7;  end
            64'b00000001????????????????????????????????????????????????????????: begin out = 10'd7;  len = 6'd8;  end
            64'b000000001???????????????????????????????????????????????????????: begin out = 10'd8;  len = 6'd9;  end
            64'b0000000001??????????????????????????????????????????????????????: begin out = 10'd9;  len = 6'd10; end
            64'b00000000001?????????????????????????????????????????????????????: begin out = 10'd10; len = 6'd11; end
            64'b000000000001????????????????????????????????????????????????????: begin out = 10'd11; len = 6'd12; end
            64'b0000000000001???????????????????????????????????????????????????: begin out = 10'd12; len = 6'd13; end
            64'b00000000000001??????????????????????????????????????????????????: begin out = 10'd13; len = 6'd14; end
            64'b000000000000001?????????????????????????????????????????????????: begin out = 10'd14; len = 6'd15; end
            64'b0000000000000001????????????????????????????????????????????????: begin out = 10'd15; len = 6'd16; end
            64'b00000000000000001???????????????????????????????????????????????: begin out = 10'd16; len = 6'd17; end
            64'b000000000000000001??????????????????????????????????????????????: begin out = 10'd17; len = 6'd18; end
            64'b0000000000000000001?????????????????????????????????????????????: begin out = 10'd18; len = 6'd19; end
            64'b00000000000000000001????????????????????????????????????????????: begin out = 10'd19; len = 6'd20; end
            64'b000000000000000000001???????????????????????????????????????????: begin out = 10'd20; len = 6'd21; end
            64'b0000000000000000000001??????????????????????????????????????????: begin out = 10'd21; len = 6'd22; end
            64'b00000000000000000000001?????????????????????????????????????????: begin out = 10'd22; len = 6'd23; end
            64'b000000000000000000000001????????????????????????????????????????: begin out = 10'd23; len = 6'd24; end
            64'b0000000000000000000000001???????????????????????????????????????: begin out = 10'd24; len = 6'd25; end
            64'b00000000000000000000000001??????????????????????????????????????: begin out = 10'd25; len = 6'd26; end
            64'b000000000000000000000000001?????????????????????????????????????: begin out = 10'd26; len = 6'd27; end
            64'b0000000000000000000000000001????????????????????????????????????: begin out = 10'd27; len = 6'd28; end
            64'b00000000000000000000000000001???????????????????????????????????: begin out = 10'd28; len = 6'd29; end
            64'b000000000000000000000000000001??????????????????????????????????: begin out = 10'd29; len = 6'd30; end
            64'b0000000000000000000000000000001?????????????????????????????????: begin out = 10'd30; len = 6'd31; end
            64'b00000000000000000000000000000001????????????????????????????????: begin out = 10'd31; len = 6'd32; end
            64'b000000000000000000000000000000001???????????????????????????????: begin out = 10'd32; len = 6'd33; end
            64'b0000000000000000000000000000000001??????????????????????????????: begin out = 10'd33; len = 6'd34; end
            64'b00000000000000000000000000000000001?????????????????????????????: begin out = 10'd34; len = 6'd35; end
            64'b000000000000000000000000000000000001????????????????????????????: begin out = 10'd35; len = 6'd36; end
            64'b0000000000000000000000000000000000001???????????????????????????: begin out = 10'd36; len = 6'd37; end
            64'b00000000000000000000000000000000000001??????????????????????????: begin out = 10'd37; len = 6'd38; end
            64'b000000000000000000000000000000000000001?????????????????????????: begin out = 10'd38; len = 6'd39; end
            64'b0000000000000000000000000000000000000001????????????????????????: begin out = 10'd39; len = 6'd40; end
            64'b00000000000000000000000000000000000000001???????????????????????: begin out = 10'd40; len = 6'd41; end
            64'b000000000000000000000000000000000000000001??????????????????????: begin out = 10'd41; len = 6'd42; end
            64'b0000000000000000000000000000000000000000001?????????????????????: begin out = 10'd42; len = 6'd43; end
            64'b00000000000000000000000000000000000000000001????????????????????: begin out = 10'd43; len = 6'd44; end
            64'b000000000000000000000000000000000000000000001???????????????????: begin out = 10'd44; len = 6'd45; end
            64'b0000000000000000000000000000000000000000000001??????????????????: begin out = 10'd45; len = 6'd46; end
            64'b00000000000000000000000000000000000000000000001?????????????????: begin out = 10'd46; len = 6'd47; end
            64'b000000000000000000000000000000000000000000000001????????????????: begin out = 10'd47; len = 6'd48; end
            64'b0000000000000000000000000000000000000000000000001???????????????: begin out = 10'd48; len = 6'd49; end
            64'b00000000000000000000000000000000000000000000000001??????????????: begin out = 10'd49; len = 6'd50; end
            64'b000000000000000000000000000000000000000000000000001?????????????: begin out = 10'd50; len = 6'd51; end
            64'b0000000000000000000000000000000000000000000000000001????????????: begin out = 10'd51; len = 6'd52; end
            64'b00000000000000000000000000000000000000000000000000001???????????: begin out = 10'd52; len = 6'd53; end
            64'b000000000000000000000000000000000000000000000000000001??????????: begin out = 10'd53; len = 6'd54; end
            64'b0000000000000000000000000000000000000000000000000000001?????????: begin out = 10'd54; len = 6'd55; end
            64'b00000000000000000000000000000000000000000000000000000001????????: begin out = 10'd55; len = 6'd56; end
            64'b000000000000000000000000000000000000000000000000000000001???????: begin out = 10'd56; len = 6'd57; end
            64'b0000000000000000000000000000000000000000000000000000000001??????: begin out = 10'd57; len = 6'd58; end
            64'b00000000000000000000000000000000000000000000000000000000001?????: begin out = 10'd58; len = 6'd59; end
            64'b000000000000000000000000000000000000000000000000000000000001????: begin out = 10'd59; len = 6'd60; end
            64'b0000000000000000000000000000000000000000000000000000000000001???: begin out = 10'd60; len = 6'd61; end
            64'b00000000000000000000000000000000000000000000000000000000000001??: begin out = 10'd61; len = 6'd62; end
            64'b000000000000000000000000000000000000000000000000000000000000001?: begin out = 10'd62; len = 6'd63; end
            64'b0000000000000000000000000000000000000000000000000000000000000001: begin out = 10'd63; len = 6'd63; end
            default: begin out = 10'd63; len = 6'd0; end
        endcase
    end
    else begin
        out <= 10'd63;
        len <= 6'd0;
    end
end

endmodule
